`define MINIMAL_FRAME_DURATION_CLKS 6661
`define MAXIMAL_STATE_DURATION_CLKS_BITS 22  